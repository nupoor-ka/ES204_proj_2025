module TestBench;
    reg [31:0] a, b;
    wire [31:0] product;
    
    fp32 uut (
        .a(a),
        .b(b),
        .product(product)
    );
    
    initial begin
        $monitor("A: %b, B: %b, Product: %d", a, b, product);
        
        a = 32'b01000000010110011001100110011010; // 3.4 in IEEE 754
        b = 32'b01000000000011001100110011001101; // 2.2 in IEEE 754
        #10;
        // product= 7.48
        a = 32'b11000000101000000000000000000000; // -5.0 in IEEE 754
        b = 32'b01000000010000000000000000000000; // 3.0 in IEEE 754
        #10;
        // product= -15
        a = 32'b01000000000000000000000000000000; // 2.0 in IEEE 754
        b = 32'b01000000000000000000000000000000; // 2.0 in IEEE 754
        #10;
        // product = 4
        a = 32'b00000000000000000000000000000000; // 0.0 in IEEE 754
        b = 32'b01000000010000000000000000000000; // 3.0 in IEEE 754
        #10;
        // product= 0
        a = 32'b01111111100000000000000000000000; // infinity 
        b = 32'b01000000010000000000000000000000; // 3.0 in IEEE 754
        #10;
        // product= +infinity
        a = 32'b01111111100000000000100000000000; // NaN
        b = 32'b01000000010000000000000000000000; // 3.0 in IEEE 754
        #10;
        // product = NaN 
        $finish;
    end
endmodule
